/* bus sizes, in bits */
`define BYTESIZE        8       /* size of a byte */
`define REGADDRSIZE     5       /* size of register address */
`define OPCODESIZE      11      /* size of largest opcode */
`define ALUOPSIZE       6       /* size of alu's operation bus */
`define FLAGSIZE        4       /* number of instruction flags */
`define WORDSIZE        64      /* size of a word */
`define INSTSIZE        32      /* size of a instruction */
`define SHAMTSIZE       6       /* size of shift amount */
`define SHORTSIZE       26      /* size of the largest possible immediate */
