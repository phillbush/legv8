/* size and bits of forwarding unit control signal */
`define FORWARDSIZE  2  /* size of the forward control signal */
`define FORWARDUSE   1  /* bit specifying whether to use forwarding */
`define FORWARDSRC   0  /* bit specifying the source of the forwarding */
