/* named registers */
`define XLR     5'd30   /* return address saved by BL instructions */
`define XZR     5'd31   /* the constant zero register */
