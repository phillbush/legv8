/* memory sizes, in bytes */
`define MEMPROGSIZE     128     /* size of the program memory */
`define MEMDATASIZE     128     /* size of the data memory */
