/* size of mov's operation bus */
`define MOVOPSIZE       3

/* last two bits of ALU operation code */
`define MOVSHIFT00      'b00
`define MOVSHIFT16      'b01
`define MOVSHIFT32      'b10
`define MOVSHIFT48      'b11
