/* size of alu's operation bus */
`define ALUOPSIZE       6

/* last two bits of ALU operation code */
`define ALUOP_AND       'b00
`define ALUOP_ORR       'b01
`define ALUOP_ADD       'b10
`define ALUOP_EOR       'b11
