`timescale 1 ps / 1 ps
module testbench();
	reg rst;
	reg clk;

	datapath dut(.rst(rst), .clk(clk));

	initial
	begin
		$dumpfile("testbench.vcd");
		$dumpvars(3, testbench);
		#1000;
		$writememh("registers.dump", dut.registerfile.registers);
		$writememh("memory.dump", dut.memdata.data);
		$finish;
	end

	/* rst */
	initial
	begin
		rst = 1'b1;
		#2; rst = ~rst;
	end

	/* rst */
	initial
	begin
		clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
		#1; clk = 1'h1;
		#1; clk = 1'h0;
	end
endmodule
