/* memory sizes, in bytes */
`define MEMPROGSIZE     64      /* size of the program memory */
`define MEMDATASIZE     64      /* size of the data memory */
