/* flags */
`define FLAGSIZE        4       /* number of instruction flags */
`define NEGATIVE        3
`define ZERO            2
`define OVERFLOW        1
`define CARRY           0
